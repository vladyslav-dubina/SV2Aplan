module example;
    initial begin
        $display("Current simulation time: %0t", $time);
    end
endmodule