module main;

    typedef enum logic [1:0] {
        IDLE,
        RUNNING,
        STOPPED
    } state_t;

    state_t current_state;

    

endmodule
