module example;
    time current_time;
    initial begin
        current_time = $time;
    end
endmodule