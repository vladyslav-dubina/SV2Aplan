module main;

    typedef enum logic [1:0] {
        IDLE,
        RUNNING,
        STOPPED
    } state_t;

    
    
    initial begin
        state_t current_state;
    end

endmodule
